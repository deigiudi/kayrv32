/*
 *  BenchRV32I -- A simple RISC-V (RV32I) Processor Core
 *  Copyright (c) 2020, Alessandro Dei Giudici <alessandro.deig@live.it>
 *  
 *  A file containing definitions for decoded instruction to be performed
 *
 *  THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
 *  AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 *  IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
 *  DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
 *  FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
 *  DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
 *  SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
 *  CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
 *  OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
 *  OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.   
 *
 */

// LOADS
`define LB		10'b0000000001
`define LH		10'b0000000010
`define LBU		10'b0000000100
`define LHU		10'b0000001000
`define LW		10'b0000010000

// STORE
`define SB		10'b0000000001
`define SH		10'b0000000010
`define SW		10'b0000000100

// IMMEDIATE
`define ADDI	10'b0000000001
`define SLLI	10'b0000000010
`define SLTI	10'b0000000100
`define SLTIU	10'b0000001000
`define XORI	10'b0000010000
`define SRLI	10'b0000100000
`define SRAI	10'b0001000000
`define ORI		10'b0010000000
`define ANDI	10'b0100000000

// REGISTER
`define ADD		10'b0000000001
`define SUB		10'b0000000010
`define SLL		10'b0000000100
`define SLT		10'b0000001000
`define SLTU	10'b0000010000
`define XOR		10'b0000100000
`define SRL		10'b0001000000
`define SRA		10'b0010000000
`define OR		10'b0100000000
`define AND		10'b1000000000
// BRANCHES
`define BEQ		10'b0000000001
`define BNE		10'b0000000010
`define BLT		10'b0000000100
`define BGE		10'b0000001000
`define BLTU	10'b0000010000
`define BGEU	10'b0000100000

// MIXED
`define AUIPC	10'b0000000001
`define LUI		10'b0000000010
`define JAL		10'b0000000100
`define JALR	10'b0000001000

// SYNC
//`define FENCE		10'b
//`define FENCE.I		10'b

// ENVIRONMENT
//`define CALL			10'b
//`define EBREAK		10'b

// CONTROL STATUS REGISTER
//`define CSRRW		10'b
//`define CSRRS		10'b
//`define CSRRC		10'b
//`define CSRRWI		10'b
//`define CSRRSI		10'b
//`define CSRRCI		10'b

// NOT SUPPORTED
`define NOTSUP	10'b0000000000
